module tb_syn_prga();

// Your testbench goes here.

endmodule: tb_syn_prga
