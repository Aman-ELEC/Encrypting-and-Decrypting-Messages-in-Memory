`timescale 1 ps / 1 ps

module tb_syn_task2();


task2 dut(CLOCK_50, KEY, SW,
          HEX0, HEX1, HEX2,
          HEX3, HEX4, HEX5,
          LEDR);
// Your testbench goes here.
initial begin

// logic [7:0] memory [0:255];
// assign memory = dut.\s|altsyncram_component|auto_generated|altsyncram1|ram_block3a0 .ram_core0.ram_core0.mem;

end



endmodule: tb_syn_task2
