module tb_syn_task5();

// Your testbench goes here.

endmodule: tb_syn_task5
