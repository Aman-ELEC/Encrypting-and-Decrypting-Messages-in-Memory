module tb_syn_task3();

// Your testbench goes here.

endmodule: tb_syn_task3
