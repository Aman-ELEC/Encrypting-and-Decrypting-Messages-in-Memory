module tb_syn_arc4();

// Your testbench goes here.

endmodule: tb_syn_arc4
